`ifndef _next_pc
`define _next_pc

module next_pc(
    output [31:0] f_valP,
    input [31:0] F_valP,
    input [5:0] f_op,
    input [31:0] f_valC
);
endmodule

`endif
