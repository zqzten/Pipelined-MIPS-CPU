`ifndef _test_reg_file
`define _test_reg_file

`timescale 1ns / 1ps

`include "../src/reg_file.v"

module test_reg_file;
endmodule

`endif
