`ifndef _test_aluB
`define _test_aluB

`timescale 1ns / 1ps

`include "../src/aluB.v"

module test_aluB;
endmodule

`endif
