`ifndef _test_srcA
`define _test_srcA

`timescale 1ns / 1ps

`include "../src/srcA.v"

module srcA;
endmodule

`endif
