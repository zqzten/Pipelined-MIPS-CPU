`ifndef _test_dstM
`define _test_dstM

`timescale 1ns / 1ps

`include "../src/dstM.v"

module test_dstM;
endmodule

`endif
