`ifndef _test_M_reg
`define _test_M_reg

`timescale 1ns / 1ps

`include "../src/M_reg"

module M_reg;
endmodule

`endif
