`ifndef _dstE
`define _dstE

module dstE(
    output [4:0] d_dstE,
    input [5:0] D_op,
    input [4:0] D_rt,
    input [4:0] D_rd
);
endmodule

`endif
