`ifndef _test_D_reg
`define _test_D_reg

`timescale 1ns / 1ps

`include "../src/D_reg.v"

module test_D_reg;
endmodule

`endif
