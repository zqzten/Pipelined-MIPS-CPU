`ifndef _F_reg
`define _F_reg

module F_reg(
    output [31:0] F_valP,
    input [31:0] f_valP,
    input clk,
    input F_stall
);
endmodule

`endif
