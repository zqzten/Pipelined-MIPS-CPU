`ifndef _test_pipeline_control
`define _test_pipeline_control

`timescale 1ns / 1ps

`include "../src/pipeline_control.v"

module test_pipeline_control;
endmodule

`endif
