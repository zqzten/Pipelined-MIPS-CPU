`ifndef _dstM
`define _dstM

module dstM(
    output [4:0] d_dstM,
    input [5:0] D_op,
    input [4:0] D_rt
);
endmodule

`endif
