`ifndef _test_fwdA
`define _test_fwdA

`timescale 1ns / 1ps

`include "../src/fwdA.v"

module test_fwdA;
endmodule

`endif
