`ifndef _test_instr_mem
`define _test_instr_mem

`timescale 1ns / 1ps

`include "../src/instr_mem.v"

module test_instr_mem;
endmodule

`endif
