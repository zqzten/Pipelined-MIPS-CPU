`ifndef _test_aluA
`define _test_aluA

`timescale 1ns / 1ps

`include "../src/aluA.v"

module test_aluA;
endmodule

`endif
