`ifndef _test_E_reg
`define _test_E_reg

`timescale 1ns / 1ps

`include "../src/E_reg.v"

module test_E_reg;
endmodule

`endif
