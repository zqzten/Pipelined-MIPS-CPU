`ifndef _data_mem
`define _data_mem

module data_mem(
    output [31:0] m_valM,
    input [5:0] M_op,
    input [31:0] M_valE,
    input [31:0] M_valA
);
endmodule

`endif
