`ifndef _srcB
`define _srcB

module srcB(
    output [4:0] d_srcB,
    input [5:0] D_op,
    input [4:0] D_rt
);
endmodule

`endif
