`ifndef _test_W_reg
`define _test_W_reg

`timescale 1ns / 1ps

`include "../src/W_reg.v"

module test_W_reg;
endmodule

`endif
