`ifndef _test_fwdB
`define _test_fwdB

`timescale 1ns / 1ps

`include "../src/fwdB.v"

module test_fwdB;
endmodule

`endif
