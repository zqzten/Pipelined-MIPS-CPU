`ifndef _aluA
`define _aluA

module aluA(
    output [31:0] e_aluA,
    input [5:0] E_op,
    input [31:0] E_valC,
    input [31:0] E_valA
);
endmodule

`endif
