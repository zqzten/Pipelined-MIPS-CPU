`ifndef _test_srcB
`define _test_srcB

`timescale 1ns / 1ps

`include "../src/srcB.v"

module test_srcB;
endmodule

`endif
