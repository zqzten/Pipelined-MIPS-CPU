`ifndef _test_alufunc
`define _test_alufunc

`timescale 1ns / 1ps

`include "../src/alufunc.v"

module test_alufunc;
endmodule

`endif
