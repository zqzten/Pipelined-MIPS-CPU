`ifndef _aluB
`define _aluB

module aluB(
    output [31:0] e_aluB,
    input [5:0] E_op,
    input [31:0] E_valB
);
endmodule

`endif
