`ifndef _pipeline_control
`define _pipeline_control

module pipeline_control(
    output F_stall,
    output D_stall,
    output E_bubble,
    input [5:0] E_op,
    input [4:0] E_dstM
);
endmodule

`endif
