`ifndef _test_next_pc
`define _test_next_pc

`timescale 1ns / 1ps

`include "../src/next_pc.v"

module test_next_pc;
endmodule

`endif
