`ifndef _test_dstE
`define _test_dstE

`timescale 1ns / 1ps

`include "../src/dstE.v"

module test_dstE;
endmodule

`endif
