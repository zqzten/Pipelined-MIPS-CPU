`ifndef _srcA
`define _srcA

module srcA(
    output [4:0] d_srcA,
    input [5:0] D_op,
    input [4:0] D_rs
);
endmodule

`endif
