`ifndef _test_data_mem
`define _test_data_mem

`timescale 1ns / 1ps

`include "../src/data_mem.v"

module test_data_mem;
endmodule

`endif
