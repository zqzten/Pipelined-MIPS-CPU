`ifndef _test_F_reg
`define _test_F_reg

`timescale 1ns / 1ps

`include "../src/F_reg.v"

module test_F_reg;
endmodule

`endif
