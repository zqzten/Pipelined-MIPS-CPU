`ifndef _test_alu
`define _test_alu

`timescale 1ns / 1ps

`include "../src/aluA.v"

module test_alu;
endmodule

`endif
