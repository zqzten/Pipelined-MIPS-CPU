`ifndef _alu
`define _alu

module alu(
    output [31:0] e_valE,
    input [31:0] e_aluA,
    input [31:0] e_aluB,
    input [5:0] e_alufunc
);
endmodule

`endif
